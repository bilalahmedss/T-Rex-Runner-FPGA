module pixel_gen(pixel_x,pixel_y,clk_div1,video_on,red,blue,green,state,mover_dino,mover);
  input [9:0] pixel_x,pixel_y;
  input clk_div1;
  input video_on;
  input [2:0]state;
  input [9:0]mover_dino;
  input [9:0]mover;
  output reg [3:0] red = 0;
  output reg [3:0] blue = 0;
  output reg [3:0] green = 0;
  wire display;
  display_lose g1(pixel_x, pixel_y, display);
  wire display1;
  display_start p1(pixel_x, pixel_y, display1);

  
  localparam px = 1;
  localparam defaultWidth = 88 * px;
  localparam defaultHeight = 94 * px;
always @(posedge clk_div1) // or posedge video_on)
begin
    if ((pixel_x <= 0) || (pixel_x >= 639))
    begin
    begin
        red <= 4'h0;
        blue <= 4'h0;
        green <= 4'h0;
    end
    else
    begin
        if (state == 3'b000)
        begin  
            if (display1)
            begin
                red <= 4'hF;
                blue <= 4'hF;
                green <= 4'hF;
            end
            else
            begin
                red <= 4'h0;
                blue <= 4'h0;
                green <= 4'h0;
            end
        end

        else if (state == 3'b001) // running
        begin
    red <= video_on ? ((pixel_x >= 0) && (pixel_x <= 639) && (pixel_y >= 375) && (pixel_y <= 380) ? 4'hF : 4'h0) : 4'h0;
    blue <= video_on ? (
        ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 89 * px))
        || ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 88 * px))
        || ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 87 * px))
        || ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 86 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 85 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 84 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 83 * px))
        || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 83 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 82 * px))
        || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 82 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 81 * px))
        || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 81 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 80 * px))
        || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 80 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 79 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 78 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 77 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 76 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 75 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 74 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 73 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 72 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 71 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 70 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 69 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 68 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 67 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 66 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 65 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 64 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 63 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 62 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 61 * px))
        || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 60 * px))
        || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 59 * px))
        || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 59 * px))
        || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 58 * px))
        || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 58 * px))
        || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 57 * px))
        || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 57 * px))
        || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 56 * px))
        || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 56 * px))
        || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 55 * px))
        || ((pixel_x > 25 + 34 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 55 * px))
        || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 54 * px))
        || ((pixel_x> 25 + 34 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 54 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 7 * px) && (pixel_y == mover_dino - 53 * px))
        || ((pixel_x> 25 + 34 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 53 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 7 * px) && (pixel_y == mover_dino - 52 * px))
        || ((pixel_x> 25 + 34 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 52 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 11 * px) && (pixel_y == mover_dino - 51 * px))
        || ((pixel_x> 25 + 28 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 51 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 11 * px) && (pixel_y == mover_dino - 50 * px))
        || ((pixel_x> 25 + 28 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 50 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 11 * px) && (pixel_y == mover_dino - 49 * px))
        || ((pixel_x> 25 + 28 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 49 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 11 * px) && (pixel_y == mover_dino - 48 * px))
        || ((pixel_x> 25 + 28 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 48 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 15 * px) && (pixel_y == mover_dino - 47 * px))  
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 47 * px))
        || ((pixel_x> 25 + 64 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 47 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 15 * px) && (pixel_y == mover_dino - 46 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 46 * px))
        || ((pixel_x> 25 + 64 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 46 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 15 * px) && (pixel_y == mover_dino - 45 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 45 * px))
        || ((pixel_x> 25 + 64 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 45 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 15 * px) && (pixel_y == mover_dino - 44 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 44 * px))
        || ((pixel_x> 25 + 64 * px) && (pixel_x<= 25 + 67 * px) && (pixel_y == mover_dino - 44 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 43 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 42 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 41 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 40 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 39 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 38 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 37 * px))
        || ((pixel_x> 25 + 4 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 36 * px))
        || ((pixel_x> 25 + 8 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 35 * px))
        || ((pixel_x> 25 + 8 * px) && (pixel_x<= 25 + 59 * px) && (pixel_y == mover_dino - 34 * px))
        || ((pixel_x> 25 + 8 * px) && (pixel_x<= 25 + 55 * px) && (pixel_y == mover_dino - 33 * px))
        || ((pixel_x> 25 + 8 * px) && (pixel_x<= 25 + 55 * px) && (pixel_y == mover_dino - 32 * px))
        || ((pixel_x> 25 + 12 * px) && (pixel_x<= 25 + 55 * px) && (pixel_y == mover_dino - 31 * px))
        || ((pixel_x> 25 + 12 * px) && (pixel_x<= 25 + 55 * px) && (pixel_y == mover_dino - 30 * px))
        || ((pixel_x> 25 + 12 * px) && (pixel_x<= 25 + 55 * px) && (pixel_y == mover_dino - 29 * px))
        || ((pixel_x> 25 + 12 * px) && (pixel_x<= 25 + 55 * px) && (pixel_y == mover_dino - 28 * px))
        || ((pixel_x> 25 + 16 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 27 * px))
        || ((pixel_x> 25 + 16 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 26 * px))
        || ((pixel_x> 25 + 16 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 25 * px))
        || ((pixel_x> 25 + 16 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 24 * px))
        || ((pixel_x> 25 + 20 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 23 * px))
        || ((pixel_x> 25 + 20 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 22 * px))
        || ((pixel_x> 25 + 20 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 21 * px))
        || ((pixel_x> 25 + 20 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 20 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 35 * px) && (pixel_y == mover_dino - 19 * px))
        || ((pixel_x> 25 + 40 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 19 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 35 * px) && (pixel_y == mover_dino - 18 * px))
        || ((pixel_x> 25 + 40 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 18 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 35 * px) && (pixel_y == mover_dino - 17 * px))
        || ((pixel_x> 25 + 40 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 17 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 35 * px) && (pixel_y == mover_dino - 16 * px))
        || ((pixel_x> 25 + 40 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 16 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 15 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 15 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 14 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 14 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 13 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 13 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 12 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 12 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 27 * px) && (pixel_y == mover_dino - 11 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 11 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 27 * px) && (pixel_y == mover_dino - 10 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 10 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 27 * px) && (pixel_y == mover_dino - 9 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 9 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 27 * px) && (pixel_y == mover_dino - 8 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 47 * px) && (pixel_y == mover_dino - 8 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 7 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 7 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 6 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 6 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 5 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 5 * px))
        || ((pixel_x> 25 + 24 * px) && (pixel_x<= 25 + 31 * px) && (pixel_y == mover_dino - 4 * px))
        || ((pixel_x> 25 + 44 * px) && (pixel_x<= 25 + 51 * px) && (pixel_y == mover_dino - 4 * px))? 4'hF:4'h0 ) : 4'h0;
        green   <= video_on ? (((pixel_x > mover + 14 * px) && (pixel_x <= mover + 19 * px) && (pixel_y == 375 - 67 * px))
        || ((pixel_x > mover + 14 * px) && (pixel_x <= mover + 19 * px) && (pixel_y == 375 - 66 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 65 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 64 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 63 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 62 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 61 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 60 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 59 * px))
        || ((pixel_x > mover + 28 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 59 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 58 * px))
        || ((pixel_x > mover + 28 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 58 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 57 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 57 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 56 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 56 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 55 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 55 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 54 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 54 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 53 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 53 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 52 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 52 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 5 * px) && (pixel_y == 375 - 51 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 51 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 51 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 5 * px) && (pixel_y == 375 - 50 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 50 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 50 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 49 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 49 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 49 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 48 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 48 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 48 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 47 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 47 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 47 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 46 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 46 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 46 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 45 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 45 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 45 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 44 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 44 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 44 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 43 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 43 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 43 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 42 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 42 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 42 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 41 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 41 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 41 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 40 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 40 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 40 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 39 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 39 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 39 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 38 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 38 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 38 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 37 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 37 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 36 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 36 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 35 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 35 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 34 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 34 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 33 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 27 * px) && (pixel_y == 375 - 33 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 32 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 27 * px) && (pixel_y == 375 - 32 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 31 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 31 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 30 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 30 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 29 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 28 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 27 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 26 * px))
        || ((pixel_x > mover + 6 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 25 * px))
        || ((pixel_x > mover + 6 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 24 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 23 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 22 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 21 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 20 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 19 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 18 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 17 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 16 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 15 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 14 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 13 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 12 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 11 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 10 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 9 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 8 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 7 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 6 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 5 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 4 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 3 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 2 * px))? 4'hF:4'h0 ) : 4'h0;
        end
        ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
        
        else if(state==3'b010) // move up
        begin  
        red   <= video_on ? ((pixel_x>=0) && (pixel_x <= 639) && ( pixel_y>=375) && (pixel_y <= 380)? 4'hF:4'h0 ) : 4'h0;
        blue   <= video_on ? (
        ((pixel_x>25+48*px)&&(pixel_x<=25+79*px)&&(pixel_y==mover_dino-89*px))
        || ((pixel_x>25+48*px)&&(pixel_x<=25+79*px)&&(pixel_y==mover_dino-88*px))
        || ((pixel_x>25+48*px)&&(pixel_x<=25+79*px)&&(pixel_y==mover_dino-87*px))
        || ((pixel_x>25+48*px)&&(pixel_x<=25+79*px)&&(pixel_y==mover_dino-86*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-85*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-84*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-83*px))
        || ((pixel_x>25+56*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-83*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-82*px))
        || ((pixel_x>25+56*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-82*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-81*px))
        || ((pixel_x>25+56*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-81*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-80*px))
        || ((pixel_x>25+56*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-80*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-79*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-78*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-77*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-76*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-75*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-74*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-73*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-72*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-71*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-70*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-69*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+83*px)&&(pixel_y==mover_dino-68*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+63*px)&&(pixel_y==mover_dino-67*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+63*px)&&(pixel_y==mover_dino-66*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+63*px)&&(pixel_y==mover_dino-65*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+63*px)&&(pixel_y==mover_dino-64*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+75*px)&&(pixel_y==mover_dino-63*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+75*px)&&(pixel_y==mover_dino-62*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+75*px)&&(pixel_y==mover_dino-61*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+75*px)&&(pixel_y==mover_dino-60*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-59*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-59*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-58*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-58*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-57*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-57*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-56*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-56*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-55*px))
        || ((pixel_x>25+34*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-55*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-54*px))
        || ((pixel_x>25+34*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-54*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-53*px))
        || ((pixel_x>25+34*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-53*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+7*px)&&(pixel_y==mover_dino-52*px))
        || ((pixel_x>25+34*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-52*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+11*px)&&(pixel_y==mover_dino-51*px))
        || ((pixel_x>25+28*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-51*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+11*px)&&(pixel_y==mover_dino-50*px))
        || ((pixel_x>25+28*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-50*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+11*px)&&(pixel_y==mover_dino-49*px))
        || ((pixel_x>25+28*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-49*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+11*px)&&(pixel_y==mover_dino-48*px))
        || ((pixel_x>25+28*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-48*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+15*px)&&(pixel_y==mover_dino-47*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-47*px))
        || ((pixel_x>25+64*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-47*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+15*px)&&(pixel_y==mover_dino-46*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-46*px))
        || ((pixel_x>25+64*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-46*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+15*px)&&(pixel_y==mover_dino-45*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-45*px))
        || ((pixel_x>25+64*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-45*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+15*px)&&(pixel_y==mover_dino-44*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-44*px))
        || ((pixel_x>25+64*px)&&(pixel_x<=25+67*px)&&(pixel_y==mover_dino-44*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-43*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-42*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-41*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-40*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-39*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-38*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-37*px))
        || ((pixel_x>25+4*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-36*px))
        || ((pixel_x>25+8*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-35*px))
        || ((pixel_x>25+8*px)&&(pixel_x<=25+59*px)&&(pixel_y==mover_dino-34*px))
        || ((pixel_x>25+8*px)&&(pixel_x<=25+55*px)&&(pixel_y==mover_dino-33*px))
        || ((pixel_x>25+8*px)&&(pixel_x<=25+55*px)&&(pixel_y==mover_dino-32*px))
        || ((pixel_x>25+12*px)&&(pixel_x<=25+55*px)&&(pixel_y==mover_dino-31*px))
        || ((pixel_x>25+12*px)&&(pixel_x<=25+55*px)&&(pixel_y==mover_dino-30*px))
        || ((pixel_x>25+12*px)&&(pixel_x<=25+55*px)&&(pixel_y==mover_dino-29*px))
        || ((pixel_x>25+12*px)&&(pixel_x<=25+55*px)&&(pixel_y==mover_dino-28*px))
        || ((pixel_x>25+16*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-27*px))
        || ((pixel_x>25+16*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-26*px))
        || ((pixel_x>25+16*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-25*px))
        || ((pixel_x>25+16*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-24*px))
        || ((pixel_x>25+20*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-23*px))
        || ((pixel_x>25+20*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-22*px))
        || ((pixel_x>25+20*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-21*px))
        || ((pixel_x>25+20*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-20*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+35*px)&&(pixel_y==mover_dino-19*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-19*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+35*px)&&(pixel_y==mover_dino-18*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-18*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+35*px)&&(pixel_y==mover_dino-17*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-17*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+35*px)&&(pixel_y==mover_dino-16*px))
        || ((pixel_x>25+40*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-16*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-15*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-15*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-14*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-14*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-13*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-13*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-12*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-12*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+27*px)&&(pixel_y==mover_dino-11*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-11*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+27*px)&&(pixel_y==mover_dino-10*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-10*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+27*px)&&(pixel_y==mover_dino-9*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-9*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+27*px)&&(pixel_y==mover_dino-8*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+47*px)&&(pixel_y==mover_dino-8*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-7*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-7*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-6*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-6*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-5*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-5*px))
        || ((pixel_x>25+24*px)&&(pixel_x<=25+31*px)&&(pixel_y==mover_dino-4*px))
        || ((pixel_x>25+44*px)&&(pixel_x<=25+51*px)&&(pixel_y==mover_dino-4*px))? 4'hF:4'h0 ) : 4'h0;
        green   <= video_on ? (((pixel_x > mover + 14 * px) && (pixel_x <= mover + 19 * px) && (pixel_y == 375 - 67 * px))
        || ((pixel_x > mover + 14 * px) && (pixel_x <= mover + 19 * px) && (pixel_y == 375 - 66 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 65 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 64 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 63 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 62 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 61 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 60 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 59 * px))
        || ((pixel_x > mover + 28 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 59 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 58 * px))
        || ((pixel_x > mover + 28 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 58 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 57 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 57 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 56 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 56 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 55 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 55 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 54 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 54 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 53 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 53 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 52 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 52 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 5 * px) && (pixel_y == 375 - 51 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 51 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 51 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 5 * px) && (pixel_y == 375 - 50 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 50 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 50 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 49 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 49 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 49 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 48 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 48 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 48 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 47 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 47 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 47 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 46 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 46 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 46 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 45 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 45 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 45 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 44 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 44 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 44 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 43 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 43 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 43 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 42 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 42 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 42 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 41 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 41 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 41 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 40 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 40 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 40 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 39 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 39 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 39 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 38 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 38 * px))
        || ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 38 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 37 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 37 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 36 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 36 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 35 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 35 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 34 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 34 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 33 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 27 * px) && (pixel_y == 375 - 33 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 32 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 27 * px) && (pixel_y == 375 - 32 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 31 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 31 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 30 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 30 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 29 * px))
        || ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 28 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 27 * px))
        || ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 26 * px))
        || ((pixel_x > mover + 6 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 25 * px))
        || ((pixel_x > mover + 6 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 24 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 23 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 22 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 21 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 20 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 19 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 18 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 17 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 16 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 15 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 14 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 13 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 12 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 11 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 10 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 9 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 8 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 7 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 6 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 5 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 4 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 3 * px))
        || ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 2 * px))? 4'hF:4'h0 ) : 4'h0;
        end
        ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
        else if(state==3'b011) //move down
        begin  
        red   <= video_on ? ((pixel_x>=0) && (pixel_x <= 639) && ( pixel_y>=375) && (pixel_y <= 380)? 4'hF:4'h0 ) : 4'h0;
        blue   <= video_on ? (
 
    ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 89 * px))
    || ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 88 * px))
    || ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 87 * px))
    || ((pixel_x > 25 + 48 * px) && (pixel_x <= 25 + 79 * px) && (pixel_y == mover_dino - 86 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 85 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 84 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 83 * px))
    || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 83 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 82 * px))
    || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 82 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 81 * px))
    || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 81 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 80 * px))
    || ((pixel_x > 25 + 56 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 80 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 79 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 78 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 77 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 76 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 75 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 74 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 73 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 72 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 71 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 70 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 69 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 83 * px) && (pixel_y == mover_dino - 68 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 67 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 66 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 65 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 63 * px) && (pixel_y == mover_dino - 64 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 63 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 62 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 61 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 75 * px) && (pixel_y == mover_dino - 60 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 59 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 59 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 58 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 58 * px))
	|| ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 57 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 57 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 56 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 56 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 55 * px))
    || ((pixel_x > 25 + 34 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 55 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 54 * px))
    || ((pixel_x > 25 + 34 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 54 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 53 * px))
    || ((pixel_x > 25 + 34 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 53 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 7 * px) && (pixel_y == mover_dino - 52 * px))
    || ((pixel_x > 25 + 34 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 52 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 11 * px) && (pixel_y == mover_dino - 51 * px))
    || ((pixel_x > 25 + 28 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 51 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 11 * px) && (pixel_y == mover_dino - 50 * px))
    || ((pixel_x > 25 + 28 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 50 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 11 * px) && (pixel_y == mover_dino - 49 * px))
    || ((pixel_x > 25 + 28 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 49 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 11 * px) && (pixel_y == mover_dino - 48 * px))
    || ((pixel_x > 25 + 28 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 48 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 15 * px) && (pixel_y == mover_dino - 47 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 47 * px))
    || ((pixel_x > 25 + 64 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 47 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 15 * px) && (pixel_y == mover_dino - 46 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 46 * px))
    || ((pixel_x > 25 + 64 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 46 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 15 * px) && (pixel_y == mover_dino - 45 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 45 * px))
    || ((pixel_x > 25 + 64 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 45 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 15 * px) && (pixel_y == mover_dino - 44 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 44 * px))
    || ((pixel_x > 25 + 64 * px) && (pixel_x <= 25 + 67 * px) && (pixel_y == mover_dino - 44 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 43 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 42 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 41 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 40 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 39 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 38 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 37 * px))
    || ((pixel_x > 25 + 4 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 36 * px))
    || ((pixel_x > 25 + 8 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 35 * px))
    || ((pixel_x > 25 + 8 * px) && (pixel_x <= 25 + 59 * px) && (pixel_y == mover_dino - 34 * px))
    || ((pixel_x > 25 + 8 * px) && (pixel_x <= 25 + 55 * px) && (pixel_y == mover_dino - 33 * px))
    || ((pixel_x > 25 + 8 * px) && (pixel_x <= 25 + 55 * px) && (pixel_y == mover_dino - 32 * px))
    || ((pixel_x > 25 + 12 * px) && (pixel_x <= 25 + 55 * px) && (pixel_y == mover_dino - 31 * px))
    || ((pixel_x > 25 + 12 * px) && (pixel_x <= 25 + 55 * px) && (pixel_y == mover_dino - 30 * px))
    || ((pixel_x > 25 + 12 * px) && (pixel_x <= 25 + 55 * px) && (pixel_y == mover_dino - 29 * px))
    || ((pixel_x > 25 + 12 * px) && (pixel_x <= 25 + 55 * px) && (pixel_y == mover_dino - 28 * px))
    || ((pixel_x > 25 + 16 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 27 * px))
    || ((pixel_x > 25 + 16 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 26 * px))
    || ((pixel_x > 25 + 16 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 25 * px))
    || ((pixel_x > 25 + 16 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 24 * px))
    || ((pixel_x > 25 + 20 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 23 * px))
    || ((pixel_x > 25 + 20 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 22 * px))
    || ((pixel_x > 25 + 20 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 21 * px))
    || ((pixel_x > 25 + 20 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 20 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 35 * px) && (pixel_y == mover_dino - 19 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 19 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 35 * px) && (pixel_y == mover_dino - 18 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 18 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 35 * px) && (pixel_y == mover_dino - 17 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 17 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 35 * px) && (pixel_y == mover_dino - 16 * px))
    || ((pixel_x > 25 + 40 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 16 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 15 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 15 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 14 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 14 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 13 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 13 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 12 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 12 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 27 * px) && (pixel_y == mover_dino - 11 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 11 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 27 * px) && (pixel_y == mover_dino - 10 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 10 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 27 * px) && (pixel_y == mover_dino - 9 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 9 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 27 * px) && (pixel_y == mover_dino - 8 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 47 * px) && (pixel_y == mover_dino - 8 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 7 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 7 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 6 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 6 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 5 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 5 * px))
    || ((pixel_x > 25 + 24 * px) && (pixel_x <= 25 + 31 * px) && (pixel_y == mover_dino - 4 * px))
    || ((pixel_x > 25 + 44 * px) && (pixel_x <= 25 + 51 * px) && (pixel_y == mover_dino - 4 * px))



 ? 4'hF:4'h0 ) : 4'h0;
        green   <= video_on ? (((pixel_x > mover + 14 * px) && (pixel_x <= mover + 19 * px) && (pixel_y == 375 - 67 * px))
	|| ((pixel_x > mover + 14 * px) && (pixel_x <= mover + 19 * px) && (pixel_y == 375 - 66 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 65 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 64 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 63 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 62 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 61 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 60 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 59 * px))
	|| ((pixel_x > mover + 28 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 59 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 58 * px))
	|| ((pixel_x > mover + 28 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 58 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 57 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 57 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 56 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 56 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 55 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 55 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 54 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 54 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 53 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 53 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 52 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 52 * px))
	|| ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 5 * px) && (pixel_y == 375 - 51 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 51 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 51 * px))
	|| ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 5 * px) && (pixel_y == 375 - 50 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 50 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 50 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 49 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 49 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 49 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 48 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 48 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 48 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 47 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 47 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 47 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 46 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 46 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 46 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 45 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 45 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 45 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 44 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 44 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 44 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 43 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 43 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 43 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 42 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 42 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 42 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 41 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 41 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 41 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 40 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 40 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 40 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 39 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 39 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 39 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 38 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 38 * px))
	|| ((pixel_x > mover + 26 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 38 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 37 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 37 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 36 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 31 * px) && (pixel_y == 375 - 36 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 35 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 35 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 34 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 29 * px) && (pixel_y == 375 - 34 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 33 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 27 * px) && (pixel_y == 375 - 33 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 32 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 27 * px) && (pixel_y == 375 - 32 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 31 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 31 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 7 * px) && (pixel_y == 375 - 30 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 30 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 29 * px))
	|| ((pixel_x > mover + 2 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 28 * px))
	|| ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 27 * px))
	|| ((pixel_x > mover + 4 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 26 * px))
	|| ((pixel_x > mover + 6 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 25 * px))
	|| ((pixel_x > mover + 6 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 24 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 23 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 22 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 21 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 20 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 19 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 18 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 17 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 16 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 15 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 14 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 13 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 12 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 11 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 10 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 9 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 8 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 7 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 6 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 5 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 4 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 3 * px))
	|| ((pixel_x > mover + 12 * px) && (pixel_x <= mover + 21 * px) && (pixel_y == 375 - 2 * px))? 4'hF:4'h0 ) : 4'h0;
        end
        else if(state==3'b100)
        begin  
         if (display) 
         begin
         red<=4'hF;
         blue<=4'hF;
         green<=4'hF;
         end
         
        
         else
         begin
         red<=4'h0;
         blue<=4'h0;
         green<=4'h0;
         end
         end
         ///////////////////////////////////
 else
 begin
 blue<=4'hF;
 end
      end
end
endmodule